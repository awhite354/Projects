magic
tech sky130A
timestamp 1644516095
<< nwell >>
rect 190 9 448 194
<< nmos >>
rect 310 -105 325 -63
<< pmos >>
rect 310 30 325 114
<< ndiff >>
rect 270 -75 310 -63
rect 270 -95 275 -75
rect 295 -95 310 -75
rect 270 -105 310 -95
rect 325 -75 360 -63
rect 325 -95 335 -75
rect 355 -95 360 -75
rect 325 -105 360 -95
<< pdiff >>
rect 270 90 310 114
rect 270 70 275 90
rect 295 70 310 90
rect 270 30 310 70
rect 325 90 360 114
rect 325 70 335 90
rect 355 70 360 90
rect 325 30 360 70
<< ndiffc >>
rect 275 -95 295 -75
rect 335 -95 355 -75
<< pdiffc >>
rect 275 70 295 90
rect 335 70 355 90
<< psubdiff >>
rect 233 -137 408 -132
rect 233 -156 270 -137
rect 290 -156 408 -137
rect 233 -162 408 -156
<< nsubdiff >>
rect 235 161 395 172
rect 235 144 265 161
rect 289 144 395 161
rect 235 141 395 144
<< psubdiffcont >>
rect 270 -156 290 -137
<< nsubdiffcont >>
rect 265 144 289 161
<< poly >>
rect 310 114 325 127
rect 310 0 325 30
rect 270 -10 325 0
rect 270 -30 280 -10
rect 300 -30 325 -10
rect 270 -40 325 -30
rect 310 -63 325 -40
rect 310 -120 325 -105
<< polycont >>
rect 280 -30 300 -10
<< locali >>
rect 264 166 294 171
rect 235 161 395 166
rect 235 160 265 161
rect 235 140 240 160
rect 260 144 265 160
rect 289 160 395 161
rect 289 144 310 160
rect 260 140 310 144
rect 330 140 370 160
rect 390 140 395 160
rect 235 136 395 140
rect 270 90 300 136
rect 270 70 275 90
rect 295 70 300 90
rect 270 30 300 70
rect 330 90 360 114
rect 330 70 335 90
rect 355 70 360 90
rect 270 -10 310 0
rect 270 -30 280 -10
rect 300 -30 310 -10
rect 270 -40 310 -30
rect 270 -75 300 -63
rect 270 -95 275 -75
rect 295 -95 300 -75
rect 270 -127 300 -95
rect 330 -75 360 70
rect 330 -95 335 -75
rect 355 -95 360 -75
rect 330 -105 360 -95
rect 233 -135 408 -127
rect 233 -155 240 -135
rect 260 -137 310 -135
rect 260 -155 270 -137
rect 233 -156 270 -155
rect 290 -155 310 -137
rect 330 -155 380 -135
rect 400 -155 408 -135
rect 290 -156 408 -155
rect 233 -162 408 -156
<< viali >>
rect 240 140 260 160
rect 310 140 330 160
rect 370 140 390 160
rect 240 -155 260 -135
rect 310 -155 330 -135
rect 380 -155 400 -135
<< metal1 >>
rect 230 160 400 170
rect 230 140 240 160
rect 260 140 310 160
rect 330 140 370 160
rect 390 140 400 160
rect 230 130 400 140
rect 230 -135 410 -125
rect 230 -155 240 -135
rect 260 -155 310 -135
rect 330 -155 380 -135
rect 400 -155 410 -135
rect 230 -165 410 -155
<< labels >>
rlabel viali 240 140 260 160 1 VDD
port 3 n
rlabel locali 270 -40 310 0 1 A
port 1 n
rlabel locali 335 -40 360 0 1 Z
port 2 n
rlabel psubdiff 238 -156 263 -133 1 GND
port 4 n
<< end >>
