magic
tech sky130A
magscale 1 2
timestamp 1644463207
<< nwell >>
rect 1861 517 1913 569
<< locali >>
rect 2777 429 2835 570
rect 440 259 682 263
rect 440 225 626 259
rect 660 225 682 259
rect 440 215 682 225
rect 1820 215 2062 263
rect 2096 215 2338 263
rect 2372 215 2614 263
rect 2645 121 2679 128
rect 2777 0 2835 141
<< viali >>
rect 863 365 897 399
rect 1387 363 1421 398
rect 30 220 67 256
rect 205 222 239 256
rect 357 219 391 253
rect 626 225 660 259
rect 728 221 762 255
rect 1237 222 1271 256
rect 1735 223 1769 257
rect 214 86 248 120
rect 1319 88 1353 122
rect 2645 87 2679 121
<< metal1 >>
rect 188 399 913 410
rect 188 365 863 399
rect 897 365 913 399
rect 188 353 913 365
rect 1363 398 1443 410
rect 1363 363 1387 398
rect 1421 363 1443 398
rect 18 256 86 265
rect 18 220 30 256
rect 67 220 86 256
rect 18 211 86 220
rect 188 256 255 353
rect 1363 351 1443 363
rect 188 222 205 256
rect 239 222 255 256
rect 188 215 255 222
rect 340 253 406 263
rect 340 219 357 253
rect 391 219 406 253
rect 340 130 406 219
rect 609 259 673 271
rect 609 225 626 259
rect 660 225 673 259
rect 609 208 673 225
rect 716 257 1786 268
rect 716 256 1735 257
rect 716 255 1237 256
rect 716 221 728 255
rect 762 222 1237 255
rect 1271 223 1735 256
rect 1769 223 1786 257
rect 1271 222 1786 223
rect 762 221 1786 222
rect 716 210 1786 221
rect 197 120 406 130
rect 197 86 214 120
rect 248 86 406 120
rect 197 76 406 86
rect 1313 122 2694 134
rect 1313 88 1319 122
rect 1353 121 2694 122
rect 1353 88 2645 121
rect 1313 87 2645 88
rect 2679 87 2694 121
rect 1313 76 2694 87
<< via1 >>
rect 24 516 76 568
rect 116 518 168 570
rect 207 520 259 572
rect 301 522 353 574
rect 386 522 438 574
rect 482 522 534 574
rect 570 522 622 574
rect 660 520 712 572
rect 758 524 810 576
rect 852 521 904 573
rect 945 522 997 574
rect 1034 521 1086 573
rect 1129 520 1181 572
rect 1219 520 1271 572
rect 1305 520 1357 572
rect 1405 521 1457 573
rect 1497 521 1549 573
rect 1588 522 1640 574
rect 1681 518 1733 570
rect 1772 518 1824 570
rect 1861 517 1913 569
rect 1955 519 2007 571
rect 2045 518 2097 570
rect 2139 517 2191 569
rect 2232 516 2284 568
rect 2322 518 2374 570
rect 2413 517 2465 569
rect 2509 517 2561 569
rect 2600 517 2652 569
rect 2691 517 2743 569
rect 2780 516 2832 568
rect 28 -18 80 34
rect 111 -28 163 24
rect 200 -25 252 27
rect 298 -25 350 27
rect 390 -27 442 25
rect 479 -28 531 24
rect 577 -27 629 25
rect 667 -28 719 24
rect 760 -25 812 27
rect 852 -34 904 18
rect 942 -26 994 26
rect 1034 -25 1086 27
rect 1128 -26 1180 26
rect 1221 -25 1273 27
rect 1302 -32 1354 20
rect 1406 -24 1458 28
rect 1494 -27 1546 25
rect 1586 -28 1638 24
rect 1681 -34 1733 18
rect 1770 -32 1822 20
rect 1863 -29 1915 23
rect 1959 -29 2011 23
rect 2046 -32 2098 20
rect 2138 -28 2190 24
rect 2229 -27 2281 25
rect 2325 -29 2377 23
rect 2415 -29 2467 23
rect 2508 -27 2560 25
rect 2599 -33 2651 19
rect 2685 -27 2737 25
rect 2776 -26 2828 26
<< metal2 >>
rect 0 576 2852 592
rect 0 574 758 576
rect 0 572 301 574
rect 0 570 207 572
rect 0 568 116 570
rect 0 516 24 568
rect 76 518 116 568
rect 168 520 207 570
rect 259 522 301 572
rect 353 522 386 574
rect 438 522 482 574
rect 534 522 570 574
rect 622 572 758 574
rect 622 522 660 572
rect 259 520 660 522
rect 712 524 758 572
rect 810 574 2852 576
rect 810 573 945 574
rect 810 524 852 573
rect 712 521 852 524
rect 904 522 945 573
rect 997 573 1588 574
rect 997 522 1034 573
rect 904 521 1034 522
rect 1086 572 1405 573
rect 1086 521 1129 572
rect 712 520 1129 521
rect 1181 520 1219 572
rect 1271 520 1305 572
rect 1357 521 1405 572
rect 1457 521 1497 573
rect 1549 522 1588 573
rect 1640 571 2852 574
rect 1640 570 1955 571
rect 1640 522 1681 570
rect 1549 521 1681 522
rect 1357 520 1681 521
rect 168 518 1681 520
rect 1733 518 1772 570
rect 1824 569 1955 570
rect 1824 518 1861 569
rect 76 517 1861 518
rect 1913 519 1955 569
rect 2007 570 2852 571
rect 2007 519 2045 570
rect 1913 518 2045 519
rect 2097 569 2322 570
rect 2097 518 2139 569
rect 1913 517 2139 518
rect 2191 568 2322 569
rect 2191 517 2232 568
rect 76 516 2232 517
rect 2284 518 2322 568
rect 2374 569 2852 570
rect 2374 518 2413 569
rect 2284 517 2413 518
rect 2465 517 2509 569
rect 2561 517 2600 569
rect 2652 517 2691 569
rect 2743 568 2852 569
rect 2743 517 2780 568
rect 2284 516 2780 517
rect 2832 516 2852 568
rect 0 496 2852 516
rect 0 34 2852 48
rect 0 -18 28 34
rect 80 28 2852 34
rect 80 27 1406 28
rect 80 24 200 27
rect 80 -18 111 24
rect 0 -28 111 -18
rect 163 -25 200 24
rect 252 -25 298 27
rect 350 25 760 27
rect 350 -25 390 25
rect 163 -27 390 -25
rect 442 24 577 25
rect 442 -27 479 24
rect 163 -28 479 -27
rect 531 -27 577 24
rect 629 24 760 25
rect 629 -27 667 24
rect 531 -28 667 -27
rect 719 -25 760 24
rect 812 26 1034 27
rect 812 18 942 26
rect 812 -25 852 18
rect 719 -28 852 -25
rect 0 -34 852 -28
rect 904 -26 942 18
rect 994 -25 1034 26
rect 1086 26 1221 27
rect 1086 -25 1128 26
rect 994 -26 1128 -25
rect 1180 -25 1221 26
rect 1273 20 1406 27
rect 1273 -25 1302 20
rect 1180 -26 1302 -25
rect 904 -32 1302 -26
rect 1354 -24 1406 20
rect 1458 26 2852 28
rect 1458 25 2776 26
rect 1458 -24 1494 25
rect 1354 -27 1494 -24
rect 1546 24 2229 25
rect 1546 -27 1586 24
rect 1354 -28 1586 -27
rect 1638 23 2138 24
rect 1638 20 1863 23
rect 1638 18 1770 20
rect 1638 -28 1681 18
rect 1354 -32 1681 -28
rect 904 -34 1681 -32
rect 1733 -32 1770 18
rect 1822 -29 1863 20
rect 1915 -29 1959 23
rect 2011 20 2138 23
rect 2011 -29 2046 20
rect 1822 -32 2046 -29
rect 2098 -28 2138 20
rect 2190 -27 2229 24
rect 2281 23 2508 25
rect 2281 -27 2325 23
rect 2190 -28 2325 -27
rect 2098 -29 2325 -28
rect 2377 -29 2415 23
rect 2467 -27 2508 23
rect 2560 19 2685 25
rect 2560 -27 2599 19
rect 2467 -29 2599 -27
rect 2098 -32 2599 -29
rect 1733 -33 2599 -32
rect 2651 -27 2685 19
rect 2737 -26 2776 25
rect 2828 -26 2852 26
rect 2737 -27 2852 -26
rect 2651 -33 2852 -27
rect 1733 -34 2852 -33
rect 0 -48 2852 -34
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636480180
transform 1 0 2760 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636480180
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636480180
transform 1 0 276 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1636480180
transform 1 0 552 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sky130_fd_sc_hd__mux2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636480180
transform 1 0 828 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1636480180
transform 1 0 1656 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1636480180
transform 1 0 1932 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1636480180
transform 1 0 2208 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1636480180
transform 1 0 2484 0 1 0
box -38 -48 314 592
<< labels >>
rlabel metal2 2 -46 2850 46 1 VGND
port 4 n
rlabel metal2 2 498 2850 590 1 VDD
port 3 n
rlabel metal1 1382 359 1429 401 1 SEL
port 2 n
rlabel metal1 22 213 83 263 1 EN
port 1 n
rlabel metal1 616 215 665 263 1 OUT
port 5 n
<< end >>
