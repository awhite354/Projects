magic
tech sky130A
timestamp 1643083951
<< nwell >>
rect 250 10 380 140
<< nmos >>
rect 310 -105 325 -63
<< pmos >>
rect 310 30 325 114
<< ndiff >>
rect 270 -75 310 -63
rect 270 -95 275 -75
rect 295 -95 310 -75
rect 270 -105 310 -95
rect 325 -75 360 -63
rect 325 -95 335 -75
rect 355 -95 360 -75
rect 325 -105 360 -95
<< pdiff >>
rect 270 90 310 114
rect 270 70 275 90
rect 295 70 310 90
rect 270 30 310 70
rect 325 90 360 114
rect 325 70 335 90
rect 355 70 360 90
rect 325 30 360 70
<< ndiffc >>
rect 275 -95 295 -75
rect 335 -95 355 -75
<< pdiffc >>
rect 275 70 295 90
rect 335 70 355 90
<< poly >>
rect 310 114 325 127
rect 310 0 325 30
rect 270 -10 325 0
rect 270 -30 280 -10
rect 300 -30 325 -10
rect 270 -40 325 -30
rect 310 -63 325 -40
rect 310 -120 325 -105
<< polycont >>
rect 280 -30 300 -10
<< locali >>
rect 260 140 310 160
rect 330 140 370 160
rect 270 90 300 140
rect 270 70 275 90
rect 295 70 300 90
rect 270 30 300 70
rect 330 90 360 114
rect 330 70 335 90
rect 355 70 360 90
rect 270 -10 310 0
rect 270 -30 280 -10
rect 300 -30 310 -10
rect 270 -40 310 -30
rect 270 -75 300 -63
rect 270 -95 275 -75
rect 295 -95 300 -75
rect 270 -135 300 -95
rect 330 -75 360 70
rect 330 -95 335 -75
rect 355 -95 360 -75
rect 330 -105 360 -95
rect 260 -155 310 -135
rect 330 -155 380 -135
<< viali >>
rect 240 140 260 160
rect 310 140 330 160
rect 370 140 390 160
rect 240 -155 260 -135
rect 310 -155 330 -135
rect 380 -155 400 -135
<< metal1 >>
rect 230 160 400 170
rect 230 140 240 160
rect 260 140 310 160
rect 330 140 370 160
rect 390 140 400 160
rect 230 130 400 140
rect 230 -135 410 -125
rect 230 -155 240 -135
rect 260 -155 310 -135
rect 330 -155 380 -135
rect 400 -155 410 -135
rect 230 -165 410 -155
<< labels >>
rlabel viali 240 -155 260 -135 1 VGND
rlabel viali 240 140 260 160 1 VDD
rlabel locali 270 -40 310 0 1 A
rlabel locali 335 -40 360 0 1 Z
<< end >>
