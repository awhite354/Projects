magic
tech sky130A
magscale 1 2
timestamp 1647376948
<< nwell >>
rect -100 -217 400 130
<< pwell >>
rect -100 -630 400 -270
<< nmos >>
rect -32 -432 -2 -304
rect 306 -432 336 -304
rect 13 -530 97 -500
rect 207 -530 291 -500
<< pmos >>
rect 13 0 97 30
rect 207 0 291 30
<< ndiff >>
rect -88 -322 -32 -304
rect -88 -356 -77 -322
rect -43 -356 -32 -322
rect -88 -432 -32 -356
rect -2 -319 97 -304
rect -2 -353 35 -319
rect 69 -353 97 -319
rect -2 -432 97 -353
rect 13 -500 97 -432
rect 207 -319 306 -304
rect 207 -353 235 -319
rect 269 -353 306 -319
rect 207 -432 306 -353
rect 336 -322 392 -304
rect 336 -356 347 -322
rect 381 -356 392 -322
rect 336 -432 392 -356
rect 207 -500 291 -432
rect 13 -546 97 -530
rect 13 -580 38 -546
rect 72 -580 97 -546
rect 13 -596 97 -580
rect 207 -546 291 -530
rect 207 -580 233 -546
rect 267 -580 291 -546
rect 207 -596 291 -580
<< pdiff >>
rect 13 75 97 86
rect 13 41 34 75
rect 68 41 97 75
rect 13 30 97 41
rect 207 75 291 86
rect 207 41 236 75
rect 270 41 291 75
rect 207 30 291 41
rect 13 -11 97 0
rect 13 -45 34 -11
rect 68 -45 97 -11
rect 13 -80 97 -45
rect 207 -11 291 0
rect 207 -45 236 -11
rect 270 -45 291 -11
rect 207 -80 291 -45
<< ndiffc >>
rect -77 -356 -43 -322
rect 35 -353 69 -319
rect 235 -353 269 -319
rect 347 -356 381 -322
rect 38 -580 72 -546
rect 233 -580 267 -546
<< pdiffc >>
rect 34 41 68 75
rect 236 41 270 75
rect 34 -45 68 -11
rect 236 -45 270 -11
<< poly >>
rect -32 0 13 30
rect 97 0 123 30
rect 181 0 207 30
rect 291 0 336 30
rect -32 -219 -2 0
rect 306 -111 336 0
rect 84 -127 336 -111
rect 84 -161 100 -127
rect 134 -141 336 -127
rect 134 -161 150 -141
rect 84 -177 150 -161
rect -32 -232 220 -219
rect -32 -249 170 -232
rect -32 -304 -2 -249
rect 154 -266 170 -249
rect 204 -266 220 -232
rect 154 -285 220 -266
rect 306 -304 336 -141
rect -32 -458 -2 -432
rect 119 -450 185 -434
rect 119 -484 135 -450
rect 169 -484 185 -450
rect 119 -500 185 -484
rect 306 -458 336 -432
rect -88 -530 13 -500
rect 97 -530 207 -500
rect 291 -530 392 -500
<< polycont >>
rect 100 -161 134 -127
rect 170 -266 204 -232
rect 135 -484 169 -450
<< locali >>
rect -60 76 364 86
rect -60 75 134 76
rect -60 41 34 75
rect 68 41 134 75
rect -60 40 134 41
rect 170 75 364 76
rect 170 41 236 75
rect 270 41 364 75
rect 170 40 364 41
rect -60 30 364 40
rect 18 -11 84 -4
rect 18 -45 34 -11
rect 68 -45 84 -11
rect 18 -111 84 -45
rect 220 -11 286 -4
rect 220 -45 236 -11
rect 270 -45 286 -11
rect 18 -127 150 -111
rect 18 -161 100 -127
rect 134 -161 150 -127
rect 18 -177 150 -161
rect -88 -322 -32 -304
rect -88 -356 -77 -322
rect -43 -356 -32 -322
rect -88 -372 -32 -356
rect 18 -319 84 -177
rect 220 -219 286 -45
rect 154 -232 286 -219
rect 154 -266 170 -232
rect 204 -266 286 -232
rect 154 -285 286 -266
rect 18 -353 35 -319
rect 69 -353 84 -319
rect 18 -400 84 -353
rect 220 -319 286 -285
rect 220 -353 235 -319
rect 269 -353 286 -319
rect 220 -400 286 -353
rect 336 -322 392 -304
rect 336 -356 347 -322
rect 381 -356 392 -322
rect 336 -372 392 -356
rect 119 -450 185 -434
rect 119 -484 135 -450
rect 169 -484 185 -450
rect 119 -500 185 -484
rect 22 -546 88 -530
rect 22 -580 38 -546
rect 72 -580 88 -546
rect 22 -596 88 -580
rect 217 -546 283 -530
rect 217 -580 233 -546
rect 267 -580 283 -546
rect 217 -596 283 -580
<< viali >>
rect 134 40 170 76
rect -77 -356 -43 -322
rect 347 -356 381 -322
rect 135 -484 169 -450
rect 38 -580 72 -546
rect 233 -580 267 -546
<< metal1 >>
rect -88 -228 -32 -218
rect -88 -280 -86 -228
rect -34 -280 -32 -228
rect -88 -322 -32 -280
rect -88 -356 -77 -322
rect -43 -356 -32 -322
rect -88 -623 -32 -356
rect 27 -546 83 86
rect 122 76 182 86
rect 122 40 134 76
rect 170 40 182 76
rect 122 30 182 40
rect 119 -441 185 -434
rect 119 -493 126 -441
rect 178 -493 185 -441
rect 119 -500 185 -493
rect 27 -580 38 -546
rect 72 -580 83 -546
rect 27 -623 83 -580
rect 221 -530 277 86
rect 336 -228 392 -218
rect 336 -280 338 -228
rect 390 -280 392 -228
rect 336 -322 392 -280
rect 336 -356 347 -322
rect 381 -356 392 -322
rect 221 -546 278 -530
rect 221 -580 233 -546
rect 267 -580 278 -546
rect 221 -623 278 -580
rect 336 -623 392 -356
<< via1 >>
rect -86 -280 -34 -228
rect 126 -450 178 -441
rect 126 -484 135 -450
rect 135 -484 169 -450
rect 169 -484 178 -450
rect 126 -493 178 -484
rect 338 -280 390 -228
<< metal2 >>
rect -88 -228 392 -218
rect -88 -280 -86 -228
rect -34 -270 338 -228
rect -34 -280 -32 -270
rect -88 -290 -32 -280
rect 336 -280 338 -270
rect 390 -280 392 -228
rect 336 -290 392 -280
rect -88 -441 392 -434
rect -88 -493 126 -441
rect 178 -493 392 -441
rect -88 -500 392 -493
<< labels >>
rlabel locali 94 -167 140 -125 1 Q
port 3 n
rlabel locali 163 -276 213 -228 1 QB
port 4 n
rlabel metal2 -84 -492 9 -445 1 WL
port 2 n
rlabel metal1 -83 -616 -39 -535 1 GND
port 1 n
rlabel metal1 341 -615 385 -534 1 GND
port 1 n
rlabel metal1 226 11 275 78 1 BR
port 6 n
rlabel metal1 30 19 78 80 1 BL
port 5 n
rlabel metal1 150 79 150 79 1 VDD
port 7 n
rlabel pwell 151 -585 151 -585 1 VNB
port 8 n
rlabel nwell 148 -41 148 -41 1 VPB
port 9 n
<< properties >>
string FIXED_BBOX -60 -623 364 58
<< end >>
